/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_Mr_Latch (
    input  wire       VGND,
    input  wire       VDPWR,    // 1.8v power supply
//    input  wire       VAPWR,    // 3.3v power supply
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    inout  wire [7:0] ua,       // Analog pins, only ua[5:0] can be used
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

wire Qn, Qn, S, R;

    assign S= ua[0];
assign R=ua[1] ;

    assign ua[2]= Q;
    assign ua[3]= Qn;

    assign ua[5:4] = 2'b00;
    //assign uo_out[7:1] = 7'b0000000; 
    assign ui_in[7:0] = 8'b00000000;


nor NOR1(Q, S, Qn);
nor NOR2(Qn, R, Q);

  //assign uio_out = 0;
    assign uio_oe  = 0;
    assign uio_in =0
  // List all unused inputs to prevent warnings
wire _unused = &{ena, clk, rst_n, 1'b0};

    
endmodule
